// Thread is a lightweight process created inside another process... sv allows multiple threads inside a single process and threads run concurrently!..
// fork... join => Start all threads in parallel and wait until every thread finishes and statement are sequentially one after another
