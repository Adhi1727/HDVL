// Array radomization
