//shallow copy
