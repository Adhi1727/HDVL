// Super keyword
