// An interface is a bundle of signals . It encapulates the signals and communication with the design and testbench components!...
