// Without super key
