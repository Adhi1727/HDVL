// base class
