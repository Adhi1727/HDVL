// we can avoid overriding
