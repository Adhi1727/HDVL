// by
