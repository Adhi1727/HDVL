//Shallow copy
